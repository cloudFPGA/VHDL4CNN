-- /*******************************************************************************
--  * Copyright 2021 -- 2024 IBM Corporation
--  *
--  * Licensed under the Apache License, Version 2.0 (the "License");
--  * you may not use this file except in compliance with the License.
--  * You may obtain a copy of the License at
--  *
--  *     http://www.apache.org/licenses/LICENSE-2.0
--  *
--  * Unless required by applicable law or agreed to in writing, software
--  * distributed under the License is distributed on an "AS IS" BASIS,
--  * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
--  * See the License for the specific language governing permissions and
--  * limitations under the License.
-- *******************************************************************************/

-- ************************************************
-- Copyright (c) 2017, Kamel ABDELOUAHAB
-- All rights reserved.
--
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions are met:
--
-- * Redistributions of source code must retain the above copyright notice, this
--   list of conditions and the following disclaimer.
--
-- * Redistributions in binary form must reproduce the above copyright notice,
--   this list of conditions and the following disclaimer in the documentation
--   and/or other materials provided with the distribution.
--
-- THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
-- AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
-- IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
-- DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE
-- FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
-- DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR
-- SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER
-- CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY,
-- OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE
-- OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- ************************************************

--  *
--  *                       VHDL4CNN
--  *    =============================================
--  *     Created/Refactored: Feb 2022
--  *     Authors: NGL
--  *     Description: Implementation of a Multiple-Constant-Multiplier:
--  *                  This IP multiplies an input array with CONSTANT
--  *                  coefficients (3D convolution kernels).
--  *

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library work;
use work.cnn_types.all;

entity MCM is
  generic(
    BITWIDTH       : integer;
    DOT_PRODUCT_SIZE : integer;
    KERNEL_VALUE     : pixel_array
    );
  port(
    clk       : in  std_logic;
    reset_n   : in  std_logic;
    enable    : in  std_logic;
    in_data   : in  pixel_array (DOT_PRODUCT_SIZE - 1 downto 0);
    in_valid  : in  std_logic;
    out_data  : out prod_array (DOT_PRODUCT_SIZE - 1 downto 0);
    out_valid : out std_logic
    );
end MCM;

architecture rtl of MCM is

begin


  process(clk)
    variable tmp_prod_result: std_logic_vector(2*BITWIDTH-1 downto 0);
  begin
    if (rising_edge(clk)) then
      --if (reset_n = '0') or (enable = '0') or (in_valid = '0') then
      --  out_data  <= (others => (others => '0'));
      --  out_valid <= '0';
      --else
        mcm_loop : for i in 0 to (DOT_PRODUCT_SIZE - 1) loop
          -- out_data(i) <= std_logic_vector(signed(KERNEL_VALUE(i)) * signed(in_data(i)));
          tmp_prod_result := std_logic_vector(signed(KERNEL_VALUE(i)) * signed(in_data(i)));
          out_data(i) <= (others => '0');
          out_data(i)(2*BITWIDTH - 2 downto 0) <= tmp_prod_result(2* BITWIDTH -2 downto 0);
          -- sign bit
          out_data(i)(out_data(i)'length-1) <= tmp_prod_result(2*BITWIDTH-1);
        end loop;
        out_valid <= in_valid;
      -- end if;
    end if;
  end process;

end architecture;

